package rvant_pkg;

/////////////////////
// Parameter Enums //
/////////////////////

typedef enum integer {
    RV32MNone = 0,
    RV32MSlow = 1,
    RV32MFast = 2
} rv32m_e;

/////////////
// Opcodes //
/////////////

typedef enum logic [6:0] {
    OPCODE_LOAD     = 7'h03,
    OPCODE_MISC_MEM = 7'h0f,
    OPCODE_OP_IMM   = 7'h13,
    OPCODE_AUIPC    = 7'h17,
    OPCODE_STORE    = 7'h23,
    OPCODE_OP       = 7'h33,
    OPCODE_LUI      = 7'h37,
    OPCODE_BRANCH   = 7'h63,
    OPCODE_JALR     = 7'h67,
    OPCODE_JAL      = 7'h6f,
    OPCODE_SYSTEM   = 7'h73
} opcode_e;

endpackage
